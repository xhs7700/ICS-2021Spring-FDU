`include "common.svh"
`include "mycpu/control.svh"
`include "mycpu/instr.svh"

module ControlUnit (
    input instr_t instr,
    input i5 branch_flag,
    output control_t control,
    output i1 ins_error
);
    control_t control_nop;
    i6 opcode,funct;
    assign opcode=instr[31:26];
    assign funct=instr[5:0];
    assign control_nop={
        ALU_SRC_NONE,
        ALU_SRC_NONE,
        ALU_OP_NONE,
        BR_NONE,
        5'b00000,
        VAL_NONE,
        REG_DST_NONE,
        LS_NONE,
        EXC_None
    };
    always_comb begin
        ins_error=1'b0;
        if (instr==32'd0) begin
            control=control_nop;
        end else begin
            control={
                ALU_SRC_RS,
                ALU_SRC_IMM_S,
                ALU_OP_NONE,
                BR_NONE,
                5'b10000,
                VAL_ALU_RES,
                REG_DST_RT,
                LS_NONE,
                EXC_None
            };
            unique case (opcode)
                OP_RTYPE: begin
                    control.alu_src_b=ALU_SRC_RT;
                    control.reg_dst=REG_DST_RD;
                    case (funct)
                        FN_ADD:begin
                            control.alu_op=ALU_OP_PLUS;
                            control.exc_flag=EXC_Ov;
                        end
                        FN_ADDU:control.alu_op=ALU_OP_PLUS;
                        FN_AND:control.alu_op=ALU_OP_AND;
                        FN_BREAK:begin
                            control.alu_src_a=ALU_SRC_NONE;
                            control.alu_src_b=ALU_SRC_NONE;
                            control.alu_op=ALU_OP_NONE;
                            control.branch=BR_NONE;
                            control.reg_write_en=1'b0;
                            control.reg_write_val=VAL_NONE;
                            control.reg_dst=REG_DST_NONE;
                            control.exc_flag=EXC_BP;
                        end
                        FN_DIV:begin
                            control.alu_op=ALU_OP_DIV;
                            control.reg_write_en=1'b0;
                            control.hilo_write_en=2'b11;
                            control.reg_write_val=VAL_MULT_RES;
                            control.reg_dst=REG_DST_NONE;
                        end
                        FN_DIVU:begin
                            control.alu_op=ALU_OP_DIVU;
                            control.reg_write_en=1'b0;
                            control.hilo_write_en=2'b11;
                            control.reg_write_val=VAL_MULT_RES;
                            control.reg_dst=REG_DST_NONE;
                        end
                        FN_JALR:begin
                            control.alu_src_b=ALU_SRC_NONE;
                            control.branch=BR_JR;
                            control.reg_write_val=VAL_PC;
                        end
                        FN_JR:begin
                            control.alu_src_b=ALU_SRC_NONE;
                            control.branch=BR_JR;
                            control.reg_write_en=1'b0;
                            control.reg_write_val=VAL_NONE;
                            control.reg_dst=REG_DST_NONE;
                        end
                        FN_MFHI:begin
                            control.alu_src_b=ALU_SRC_HI;
                            control.alu_op=ALU_OP_OR;
                        end
                        FN_MFLO:begin
                            control.alu_src_b=ALU_SRC_LO;
                            control.alu_op=ALU_OP_OR;
                        end
                        FN_MTHI:begin
                            control.alu_src_b=ALU_SRC_ZERO;
                            control.alu_op=ALU_OP_OR;
                            control.reg_write_en=1'b0;
                            control.hilo_write_en=2'b10;
                            control.reg_dst=REG_DST_NONE;
                        end
                        FN_MTLO:begin
                            control.alu_src_b=ALU_SRC_ZERO;
                            control.alu_op=ALU_OP_OR;
                            control.reg_write_en=1'b0;
                            control.hilo_write_en=2'b01;
                            control.reg_dst=REG_DST_NONE;
                        end
                        FN_MULT:begin
                            control.alu_op=ALU_OP_MULT;
                            control.reg_write_en=1'b0;
                            control.hilo_write_en=2'b11;
                            control.reg_write_val=VAL_MULT_RES;
                            control.reg_dst=REG_DST_NONE;
                        end
                        FN_MULTU:begin
                            control.alu_op=ALU_OP_MULTU;
                            control.reg_write_en=1'b0;
                            control.hilo_write_en=2'b11;
                            control.reg_write_val=VAL_MULT_RES;
                            control.reg_dst=REG_DST_NONE;
                        end
                        FN_NOR:control.alu_op=ALU_OP_NOR;
                        FN_OR:control.alu_op=ALU_OP_OR;
                        FN_SLL:begin
                            control.alu_op=ALU_OP_SLL;
                            control.alu_src_a=ALU_SRC_SHAMT;
                            control.alu_src_b=ALU_SRC_RT;
                        end
                        FN_SLLV:control.alu_op=ALU_OP_SLLV;
                        FN_SLT:control.alu_op=ALU_OP_SLT;
                        FN_SLTU:control.alu_op=ALU_OP_SLTU;
                        FN_SRA:begin
                            control.alu_op=ALU_OP_SRA;
                            control.alu_src_a=ALU_SRC_SHAMT;
                            control.alu_src_b=ALU_SRC_RT;
                        end
                        FN_SRAV:control.alu_op=ALU_OP_SRAV;
                        FN_SRL:begin
                            control.alu_op=ALU_OP_SRL;
                            control.alu_src_a=ALU_SRC_SHAMT;
                            control.alu_src_b=ALU_SRC_RT;
                        end
                        FN_SRLV:control.alu_op=ALU_OP_SRLV;
                        FN_SUB:begin
                            control.alu_op=ALU_OP_MINUS;
                            control.exc_flag=EXC_Ov;
                        end
                        FN_SUBU:control.alu_op=ALU_OP_MINUS;
                        FN_SYSCALL:begin
                            control.alu_src_a=ALU_SRC_NONE;
                            control.alu_src_b=ALU_SRC_NONE;
                            control.alu_op=ALU_OP_NONE;
                            control.branch=BR_NONE;
                            control.reg_write_en=1'b0;
                            control.reg_write_val=VAL_NONE;
                            control.reg_dst=REG_DST_NONE;
                            control.exc_flag=EXC_Sys;
                        end
                        FN_XOR:control.alu_op=ALU_OP_XOR;
                        default:begin
                            control=control_nop;
                            ins_error=1'b1;
                        end
                    endcase
                end
                OP_BTYPE: begin
                    control.alu_src_b=ALU_SRC_ZERO;
                    control.reg_write_en=1'b0;
                    control.reg_write_val=VAL_NONE;
                    control.reg_dst=REG_DST_NONE;
                    case (branch_flag)
                        BF_BGEZ:control.branch=BR_BGEZ;
                        BF_BLTZ:control.branch=BR_BLTZ;
                        BF_BGEZAL:begin
                            control.branch=BR_BGEZ;
                            control.reg_write_en=1'b1;
                            control.reg_write_val=VAL_PC;
                            control.reg_dst=REG_DST_RA;
                        end
                        BF_BLTZAL:begin
                            control.branch=BR_BLTZ;
                            control.reg_write_en=1'b1;
                            control.reg_write_val=VAL_PC;
                            control.reg_dst=REG_DST_RA;
                        end
                        default:control=control_nop;
                    endcase
                end
                OP_COP0:begin
                    case (instr[25:21])
                        control.alu_src_a=ALU_SRC_NONE;
                        5'b10000:begin // ERET
                            control.alu_src_b=ALU_SRC_NONE;
                            control.reg_write_en=1'b0;
                            control.reg_write_val=VAL_NONE;
                            control.reg_dst=REG_DST_NONE;
                            control.exc_flag=EXC_Eret;
                        end
                        5'b00000:begin // MFC0
                            control.alu_src_b=ALU_SRC_C0;
                            control.alu_op=ALU_OP_OR;
                        end
                        5'b00100:begin // MTC0
                            control.alu_src_b=ALU_SRC_RT;
                            control.alu_op=ALU_OP_OR;
                            control.reg_write_en=1'b0;
                            control.c0_write_en=1'b1;
                            control.reg_dst=REG_DST_RD;
                        end
                    endcase
                end
                OP_ADDI:begin
                    control.alu_op=ALU_OP_PLUS;
                    control.exc_flag=EXC_Ov;
                end
                OP_ADDIU:control.alu_op=ALU_OP_PLUS;
                OP_ANDI:begin
                    control.alu_src_b=ALU_SRC_IMM_Z;
                    control.alu_op=ALU_OP_AND;
                end
                OP_BEQ:begin
                    control.alu_src_b=ALU_SRC_RT;
                    control.branch=BR_BEQ;
                    control.reg_write_en=1'b0;
                    control.reg_write_val=VAL_NONE;
                    control.reg_dst=REG_DST_NONE;
                end
                OP_BGTZ:begin
                    control.alu_src_b=ALU_SRC_ZERO;
                    control.branch=BR_BGTZ;
                    control.reg_write_en=1'b0;
                    control.reg_write_val=VAL_NONE;
                    control.reg_dst=REG_DST_NONE;
                end
                OP_BLEZ:begin
                    control.alu_src_b=ALU_SRC_ZERO;
                    control.branch=BR_BLEZ;
                    control.reg_write_en=1'b0;
                    control.reg_write_val=VAL_NONE;
                    control.reg_dst=REG_DST_NONE;
                end
                OP_BNE:begin
                    control.alu_src_b=ALU_SRC_RT;
                    control.branch=BR_BNE;
                    control.reg_write_en=1'b0;
                    control.reg_write_val=VAL_NONE;
                    control.reg_dst=REG_DST_NONE;
                end
                OP_J:begin
                    control={
                        ALU_SRC_NONE,
                        ALU_SRC_NONE,
                        ALU_OP_NONE,
                        BR_J,
                        5'b00000,
                        VAL_NONE,
                        REG_DST_NONE,
                        LS_NONE,
                        EXC_None
                    };
                end
                OP_JAL:begin
                    control={
                        ALU_SRC_NONE,
                        ALU_SRC_NONE,
                        ALU_OP_NONE,
                        BR_J,
                        5'b10000,
                        VAL_PC,
                        REG_DST_RA,
                        LS_NONE,
                        EXC_None
                    };
                end
                OP_LUI:begin
                    control.alu_src_b=ALU_SRC_IMM_H;
                    control.alu_op=ALU_OP_OR;
                end
                OP_LB:begin
                    control.alu_op=ALU_OP_PLUS;
                    control.reg_write_val=VAL_MEM;
                    control.ls_flag=LS_BTYE;
                end
                OP_LBU:begin
                    control.alu_op=ALU_OP_PLUS;
                    control.reg_write_val=VAL_MEM;
                    control.ls_flag=LS_BTYE_U;
                end
                OP_LH:begin
                    control.alu_op=ALU_OP_PLUS;
                    control.reg_write_val=VAL_MEM;
                    control.ls_flag=LS_HALFW;
                end
                OP_LHU:begin
                    control.alu_op=ALU_OP_PLUS;
                    control.reg_write_val=VAL_MEM;
                    control.ls_flag=LS_HALFW_U;
                end
                OP_LW:begin
                    control.alu_op=ALU_OP_PLUS;
                    control.reg_write_val=VAL_MEM;
                    control.ls_flag=LS_WORD;
                end
                OP_ORI:begin
                    control.alu_src_b=ALU_SRC_IMM_Z;
                    control.alu_op=ALU_OP_OR;
                end
                OP_SLTI:begin
                    control.alu_op=ALU_OP_SLT;
                end
                OP_SLTIU:begin
                    control.alu_op=ALU_OP_SLTU;
                end
                OP_SB:begin
                    control.alu_op=ALU_OP_PLUS;
                    control.reg_write_en=1'b0;
                    control.mem_write_en=1'b1;
                    control.reg_write_val=VAL_NONE;
                    control.reg_dst=REG_DST_NONE;
                    control.ls_flag=LS_BTYE;
                end
                OP_SH:begin
                    control.alu_op=ALU_OP_PLUS;
                    control.reg_write_en=1'b0;
                    control.mem_write_en=1'b1;
                    control.reg_write_val=VAL_NONE;
                    control.reg_dst=REG_DST_NONE;
                    control.ls_flag=LS_HALFW;
                end
                OP_SW:begin
                    control.alu_op=ALU_OP_PLUS;
                    control.reg_write_en=1'b0;
                    control.mem_write_en=1'b1;
                    control.reg_write_val=VAL_NONE;
                    control.reg_dst=REG_DST_NONE;
                    control.ls_flag=LS_WORD;
                end
                OP_XORI:begin
                    control.alu_src_b=ALU_SRC_IMM_Z;
                    control.alu_op=ALU_OP_XOR;
                end
                default:begin
                    control=control_nop;
                    ins_error=1'b1;
                end
            endcase
        end
    end
endmodule
`include "common.svh"
`include "mycpu/control.svh"
`include "mycpu/instr.svh"

module ControlUnit (
    input opcode_t opcode,
    input funct_t funct,
    output control_t control
);
    always_comb begin
        control={
            ALU_SRC_RS,
            ALU_SRC_IMM_S,
            ALU_OP_NONE,
            BR_NONE,
            2'b10,
            VAL_ALU_RES,
            REG_DST_RT
        };
        unique case (opcode)
            OP_RTYPE: begin
                control.alu_src_b=ALU_SRC_RT;
                control.reg_dst=REG_DST_RD;
                case (funct)
                    FN_ADDU: begin
                        control.alu_op=ALU_OP_PLUS;
                    end
                    FN_AND:begin
                        control.alu_op=ALU_OP_AND;
                    end
                    FN_JR:begin
                        control={
                            ALU_SRC_RS,
                            ALU_SRC_NONE,
                            ALU_OP_NONE,
                            BR_JR,
                            2'b00,
                            VAL_NONE,
                            REG_DST_NONE
                        };
                    end
                    FN_NOR:begin
                        control.alu_op=ALU_OP_NOR;
                    end
                    FN_OR:begin
                        control.alu_op=ALU_OP_OR;
                    end
                    FN_SLL:begin
                        control.alu_op=ALU_OP_SLL;
                        control.alu_src_a=ALU_SRC_SHAMT;
                        control.alu_src_b=ALU_SRC_RT;
                    end
                    FN_SLT:begin
                        control.alu_op=ALU_OP_SLT;
                    end
                    FN_SLTU:begin
                        control.alu_op=ALU_OP_SLTU;
                    end
                    FN_SRA:begin
                        control.alu_op=ALU_OP_SRA;
                        control.alu_src_a=ALU_SRC_SHAMT;
                        control.alu_src_b=ALU_SRC_RT;
                    end
                    FN_SRL:begin
                        control.alu_op=ALU_OP_SRL;
                        control.alu_src_a=ALU_SRC_SHAMT;
                        control.alu_src_b=ALU_SRC_RT;
                    end
                    FN_SUBU:begin
                        control.alu_op=ALU_OP_MINUS;
                    end
                    FN_XOR:begin
                        control.alu_op=ALU_OP_XOR;
                    end
                    default: begin
                        control={
                            ALU_SRC_NONE,
                            ALU_SRC_NONE,
                            ALU_OP_NONE,
                            BR_NONE,
                            2'b00,
                            VAL_NONE,
                            REG_DST_NONE
                        };
                    end
                endcase
            end
            OP_ADDIU:begin
                control.alu_op=ALU_OP_PLUS;
            end
            OP_ANDI:begin
                control.alu_src_b=ALU_SRC_IMM_Z;
                control.alu_op=ALU_OP_AND;
            end
            OP_BEQ:begin
                control={
                    ALU_SRC_RS,
                    ALU_SRC_RT,
                    ALU_OP_NONE,
                    BR_BEQ,
                    2'b00,
                    VAL_NONE,
                    REG_DST_NONE
                };
            end
            OP_BNE:begin
                control={
                    ALU_SRC_RS,
                    ALU_SRC_RT,
                    ALU_OP_NONE,
                    BR_BNE,
                    2'b00,
                    VAL_NONE,
                    REG_DST_NONE
                };
            end
            OP_J:begin
                control={
                    ALU_SRC_NONE,
                    ALU_SRC_NONE,
                    ALU_OP_NONE,
                    BR_J,
                    2'b00,
                    VAL_NONE,
                    REG_DST_NONE
                };
            end
            OP_JAL:begin
                control={
                    ALU_SRC_NONE,
                    ALU_SRC_NONE,
                    ALU_OP_NONE,
                    BR_J,
                    2'b10,
                    VAL_PC,
                    REG_DST_RA
                };
            end
            OP_LUI:begin
                control.alu_src_b=ALU_SRC_IMM_H;
                control.alu_op=ALU_OP_OR;
            end
            OP_LW:begin
                control.alu_op=ALU_OP_PLUS;
                control.reg_write_val=VAL_MEM;
            end
            OP_ORI:begin
                control.alu_src_b=ALU_SRC_IMM_Z;
                control.alu_op=ALU_OP_OR;
            end
            OP_SLTI:begin
                control.alu_op=ALU_OP_SLT;
            end
            OP_SLTIU:begin
                control.alu_op=ALU_OP_SLTU;
            end
            OP_SW:begin
                control.alu_op=ALU_OP_PLUS;
                control.reg_write_en=1'b0;
                control.mem_write_en=1'b1;
                control.reg_write_val=VAL_NONE;
                control.reg_dst=REG_DST_NONE;
            end
            OP_XORI:begin
                control.alu_src_b=ALU_SRC_IMM_Z;
                control.alu_op=ALU_OP_XOR;
            end
            default: begin
                control={
                    ALU_SRC_NONE,
                    ALU_SRC_NONE,
                    ALU_OP_NONE,
                    BR_NONE,
                    2'b00,
                    VAL_NONE,
                    REG_DST_NONE
                };
            end
        endcase
    end
endmodule